library ieee;
USE ieee.std_logic_1164.all;

entity bcd7s is
port(
	bcdc:
